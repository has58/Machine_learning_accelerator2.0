Library IEEE;
use IEEE.std_logic_1164.ALL;

package My_ANN_Lib is
	
	Type integer_array is array(0 to 9) of integer;
	Type integer_matrix is array(0 to 9) of integer_array;
end package;
